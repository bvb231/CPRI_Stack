module ARP_Responder
